module controle(
    input CLK,
    input CLR,
    input [3:0] opcode,

    output reg NHLT,
    output reg HLT,
    output reg Cp,
    output reg Ep,
    output reg Lm,
    output reg CE,
    output reg L1,
    output reg Ei,
    output reg La,
    output reg Ea,
    output reg Su,
    output reg Lb,
    output reg L0
);



endmodule